module deco4_16(input [3:0] A,output logic [15:0] R);
	always@(A)
	begin case(A)
		4'd0 : R = 16'b0000000000000001;//R0
		4'd1 : R = 16'b0000000000000010;//R1
		4'd2 : R = 16'b0000000000000100;//R2
		4'd3 : R = 16'b0000000000001000;//R3
		4'd4 : R = 16'b0000000000010000;//R4
		4'd5 : R = 16'b0000000000100000;//R5
		4'd6 : R = 16'b0000000001000000;//R6
		4'd7 : R = 16'b0000000010000000;//R7
		4'd8 : R = 16'b0000000100000000;//R8
		4'd9 : R = 16'b0000001000000000;//R9
		4'd10 : R =16'b0000010000000000;//R10
		4'd11 : R =16'b0000100000000000;//R11
		4'd12 : R =16'b0001000000000000;//R12
		4'd13 : R =16'b0010000000000000;//R13
		4'd14 : R =16'b0100000000000000;//R14
		4'd15 : R =16'b1000000000000000;//R15
		default: R =16'b0000000000000000;//0
	endcase
	end
endmodule